package uart_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "uart_seq_item.sv"
	`include "uart_sequence.sv"
	`include "uart_sequencer.sv"
	`include "uart_driver.sv"
	`include "uart_agent.sv"
	`include "uart_env.sv"
	`include "uart_test.sv"
endpackage
